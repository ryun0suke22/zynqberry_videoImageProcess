module test(test_in, test_out);
input test_in;
output test_out;

assign test_out = test_in;

endmodule
